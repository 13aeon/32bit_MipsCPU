
module ROM (addr,data);
input [31:0] addr;
output reg [31:0] data;
//localparam ROM_SIZE = 32;
//reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[8:2])	//Address Must Be Word Aligned.
        0:      data <= 32'h08000003;    //0x0   j Main
        1:      data <= 32'h08000030;    //0x4   j Interrupt
        2:      data <= 32'h0800007b;    //0x8   j Exception
        3:      data <= 32'h3c164000;    //0xc   lui $s6,16384
        4:      data <= 32'h3c08ffff;    //0x10  lui $t0,65535
        5:      data <= 32'h00000000;    //0x14  sll $zero,$zero,0
        6:      data <= 32'h2108fc17;    //0x18  addi $t0,$t0,64535
        7:      data <= 32'h00000000;    //0x1c  sll $zero,$zero,0
        8:      data <= 32'h00000000;    //0x20  sll $zero,$zero,0
        9:      data <= 32'haec80000;    //0x24  sw $t0,0($s6)
        10:     data <= 32'haec80004;    //0x28  sw $t0,4($s6)
        11:     data <= 32'h20080003;    //0x2c  addi $t0,$zero,3
        12:     data <= 32'h00000000;    //0x30  sll $zero,$zero,0
        13:     data <= 32'haec80008;    //0x34  sw $t0,8($s6)
        14:     data <= 32'h20100040;    //0x38  addi $s0,$zero,64
        15:     data <= 32'hac100028;    //0x3c  sw $s0,40($zero)
        16:     data <= 32'h20100079;    //0x40  addi $s0,$zero,121
        17:     data <= 32'hac10002c;    //0x44  sw $s0,44($zero)
        18:     data <= 32'h20100024;    //0x48  addi $s0,$zero,36
        19:     data <= 32'hac100030;    //0x4c  sw $s0,48($zero)
        20:     data <= 32'h20100030;    //0x50  addi $s0,$zero,48
        21:     data <= 32'hac100034;    //0x54  sw $s0,52($zero)
        22:     data <= 32'h20100019;    //0x58  addi $s0,$zero,25
        23:     data <= 32'hac100038;    //0x5c  sw $s0,56($zero)
        24:     data <= 32'h20100012;    //0x60  addi $s0,$zero,18
        25:     data <= 32'hac10003c;    //0x64  sw $s0,60($zero)
        26:     data <= 32'h20100002;    //0x68  addi $s0,$zero,2
        27:     data <= 32'hac100040;    //0x6c  sw $s0,64($zero)
        28:     data <= 32'h20100078;    //0x70  addi $s0,$zero,120
        29:     data <= 32'hac100044;    //0x74  sw $s0,68($zero)
        30:     data <= 32'h20100000;    //0x78  addi $s0,$zero,0
        31:     data <= 32'hac100048;    //0x7c  sw $s0,72($zero)
        32:     data <= 32'h20100010;    //0x80  addi $s0,$zero,16
        33:     data <= 32'hac10004c;    //0x84  sw $s0,76($zero)
        34:     data <= 32'h20100008;    //0x88  addi $s0,$zero,8
        35:     data <= 32'hac100050;    //0x8c  sw $s0,80($zero)
        36:     data <= 32'h20100003;    //0x90  addi $s0,$zero,3
        37:     data <= 32'hac100054;    //0x94  sw $s0,84($zero)
        38:     data <= 32'h20100046;    //0x98  addi $s0,$zero,70
        39:     data <= 32'hac100058;    //0x9c  sw $s0,88($zero)
        40:     data <= 32'h20100021;    //0xa0  addi $s0,$zero,33
        41:     data <= 32'hac10005c;    //0xa4  sw $s0,92($zero)
        42:     data <= 32'h20100006;    //0xa8  addi $s0,$zero,6
        43:     data <= 32'hac100060;    //0xac  sw $s0,96($zero)
        44:     data <= 32'h2010000e;    //0xb0  addi $s0,$zero,14
        45:     data <= 32'hac100064;    //0xb4  sw $s0,100($zero)
        46:     data <= 32'h20030001;    //0xb8  addi $v1,$zero,1
        47:     data <= 32'h0800007c;    //0xbc  j End
        48:     data <= 32'h20080003;    //0xc0  addi $t0,$zero,3
        49:     data <= 32'haec80008;    //0xc4  sw $t0,8($s6)
        50:     data <= 32'h00035842;    //0xc8  srl $t3,$v1,1
        51:     data <= 32'h11600006;    //0xcc  beq $t3,$zero,A
        52:     data <= 32'h000b5842;    //0xd0  srl $t3,$t3,1
        53:     data <= 32'h1160000d;    //0xd4  beq $t3,$zero,B
        54:     data <= 32'h000b5842;    //0xd8  srl $t3,$t3,1
        55:     data <= 32'h11600014;    //0xdc  beq $t3,$zero,C
        56:     data <= 32'h000b5842;    //0xe0  srl $t3,$t3,1
        57:     data <= 32'h1160001b;    //0xe4  beq $t3,$zero,D
        58:     data <= 32'h8ecc0018;    //0xe8  lw $t4,24($s6)
        59:     data <= 32'h318c000f;    //0xec  andi $t4,$t4,15
        60:     data <= 32'h000c6080;    //0xf0  sll $t4,$t4,2
        61:     data <= 32'h8d8c0028;    //0xf4  lw $t4,40($t4)
        62:     data <= 32'h00036a00;    //0xf8  sll $t5,$v1,8
        63:     data <= 32'h01ac6020;    //0xfc  add $t4,$t5,$t4
        64:     data <= 32'haecc0014;    //0x100 sw $t4,20($s6)
        65:     data <= 32'h20030002;    //0x104 addi $v1,$zero,2
        66:     data <= 32'h0800005e;    //0x108 j cycle
        67:     data <= 32'h8ecc0018;    //0x10c lw $t4,24($s6)
        68:     data <= 32'h318c00f0;    //0x110 andi $t4,$t4,240
        69:     data <= 32'h000c6082;    //0x114 srl $t4,$t4,2
        70:     data <= 32'h8d8c0028;    //0x118 lw $t4,40($t4)
        71:     data <= 32'h00036a00;    //0x11c sll $t5,$v1,8
        72:     data <= 32'h01ac6020;    //0x120 add $t4,$t5,$t4
        73:     data <= 32'haecc0014;    //0x124 sw $t4,20($s6)
        74:     data <= 32'h20030004;    //0x128 addi $v1,$zero,4
        75:     data <= 32'h0800005e;    //0x12c j cycle
        76:     data <= 32'h8ecc001c;    //0x130 lw $t4,28($s6)
        77:     data <= 32'h318c000f;    //0x134 andi $t4,$t4,15
        78:     data <= 32'h000c6080;    //0x138 sll $t4,$t4,2
        79:     data <= 32'h8d8c0028;    //0x13c lw $t4,40($t4)
        80:     data <= 32'h00036a00;    //0x140 sll $t5,$v1,8
        81:     data <= 32'h01ac6020;    //0x144 add $t4,$t5,$t4
        82:     data <= 32'haecc0014;    //0x148 sw $t4,20($s6)
        83:     data <= 32'h20030008;    //0x14c addi $v1,$zero,8
        84:     data <= 32'h0800005e;    //0x150 j cycle
        85:     data <= 32'h8ecc001c;    //0x154 lw $t4,28($s6)
        86:     data <= 32'h318c00f0;    //0x158 andi $t4,$t4,240
        87:     data <= 32'h000c6082;    //0x15c srl $t4,$t4,2
        88:     data <= 32'h8d8c0028;    //0x160 lw $t4,40($t4)
        89:     data <= 32'h00036a00;    //0x164 sll $t5,$v1,8
        90:     data <= 32'h01ac6020;    //0x168 add $t4,$t5,$t4
        91:     data <= 32'haecc0014;    //0x16c sw $t4,20($s6)
        92:     data <= 32'h20030001;    //0x170 addi $v1,$zero,1
        93:     data <= 32'h0800005e;    //0x174 j cycle
        94:     data <= 32'h8ec80024;    //0x178 lw $t0,36($s6)
        95:     data <= 32'h00000000;    //0x17c sll $zero,$zero,0
        96:     data <= 32'h000847c0;    //0x180 sll $t0,$t0,31
        97:     data <= 32'h000847c2;    //0x184 srl $t0,$t0,31
        98:     data <= 32'h11000017;    //0x188 beq $t0,$zero,InEnd
        99:     data <= 32'h00004020;    //0x18c add $t0,$zero,$zero
        100:    data <= 32'haec80024;    //0x190 sw $t0,36($s6)
        101:    data <= 32'h8ec90018;    //0x194 lw $t1,24($s6)
        102:    data <= 32'h8eca001c;    //0x198 lw $t2,28($s6)
        103:    data <= 32'h11200008;    //0x19c beq $t1,$zero,end1
        104:    data <= 32'h11400007;    //0x1a0 beq $t2,$zero,end1
        105:    data <= 32'h112a0007;    //0x1a4 beq $t1,$t2,end2
        106:    data <= 32'h0149402a;    //0x1a8 slt $t0,$t2,$t1
        107:    data <= 32'h11000002;    //0x1ac beq $t0,$zero,loop2
        108:    data <= 32'h012a4822;    //0x1b0 sub $t1,$t1,$t2
        109:    data <= 32'h08000069;    //0x1b4 j loop1
        110:    data <= 32'h01495022;    //0x1b8 sub $t2,$t2,$t1
        111:    data <= 32'h08000069;    //0x1bc j loop1
        112:    data <= 32'h00005020;    //0x1c0 add $t2,$zero,$zero
        113:    data <= 32'h01401020;    //0x1c4 add $v0,$t2,$zero
        114:    data <= 32'haec20020;    //0x1c8 sw $v0,32($s6)
        115:    data <= 32'haec2000c;    //0x1cc sw $v0,12($s6)
        116:    data <= 32'h8ec80024;    //0x1d0 lw $t0,36($s6)
        117:    data <= 32'h00000000;    //0x1d4 sll $zero,$zero,0
        118:    data <= 32'h00084082;    //0x1d8 srl $t0,$t0,2
        119:    data <= 32'h15000002;    //0x1dc bne $t0,$zero,InEnd
        120:    data <= 32'h200a0002;    //0x1e0 addi $t2,$zero,2
        121:    data <= 32'haeca0024;    //0x1e4 sw $t2,36($s6)
        122:    data <= 32'h03400008;    //0x1e8 jr $k0
        123:    data <= 32'h03400008;    //0x1ec jr $k0
        124:    data <= 32'h0800007c;    //0x1f0 j End
      default:  data <= 32'h08000000;
    endcase
endmodule
