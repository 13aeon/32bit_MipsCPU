
module ROM (addr,data);
input [31:0] addr;
output reg [31:0] data;
//localparam ROM_SIZE = 32;
//reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[8:2])	//Address Must Be Word Aligned.
        0:      data <= 32'h08000003;    //0x0   j Main
        1:      data <= 32'h0800002c;    //0x4   j Interrupt
        2:      data <= 32'h08000076;    //0x8   j Exception
        3:      data <= 32'h3c164000;    //0xc   lui $s6,16384
        4:      data <= 32'h3c08ffff;    //0x10  lui $t0,65535
        5:      data <= 32'h2108fc17;    //0x14  addi $t0,$t0,64535
        6:      data <= 32'haec80000;    //0x18  sw $t0,0($s6)
        7:      data <= 32'haec80004;    //0x1c  sw $t0,4($s6)
        8:      data <= 32'h20080003;    //0x20  addi $t0,$zero,3
        9:      data <= 32'haec80008;    //0x24  sw $t0,8($s6)
        10:     data <= 32'h20100040;    //0x28  addi $s0,$zero,64
        11:     data <= 32'hac100028;    //0x2c  sw $s0,40($zero)
        12:     data <= 32'h20100079;    //0x30  addi $s0,$zero,121
        13:     data <= 32'hac10002c;    //0x34  sw $s0,44($zero)
        14:     data <= 32'h20100024;    //0x38  addi $s0,$zero,36
        15:     data <= 32'hac100030;    //0x3c  sw $s0,48($zero)
        16:     data <= 32'h20100030;    //0x40  addi $s0,$zero,48
        17:     data <= 32'hac100034;    //0x44  sw $s0,52($zero)
        18:     data <= 32'h20100019;    //0x48  addi $s0,$zero,25
        19:     data <= 32'hac100038;    //0x4c  sw $s0,56($zero)
        20:     data <= 32'h20100012;    //0x50  addi $s0,$zero,18
        21:     data <= 32'hac10003c;    //0x54  sw $s0,60($zero)
        22:     data <= 32'h20100002;    //0x58  addi $s0,$zero,2
        23:     data <= 32'hac100040;    //0x5c  sw $s0,64($zero)
        24:     data <= 32'h20100078;    //0x60  addi $s0,$zero,120
        25:     data <= 32'hac100044;    //0x64  sw $s0,68($zero)
        26:     data <= 32'h20100000;    //0x68  addi $s0,$zero,0
        27:     data <= 32'hac100048;    //0x6c  sw $s0,72($zero)
        28:     data <= 32'h20100010;    //0x70  addi $s0,$zero,16
        29:     data <= 32'hac10004c;    //0x74  sw $s0,76($zero)
        30:     data <= 32'h20100008;    //0x78  addi $s0,$zero,8
        31:     data <= 32'hac100050;    //0x7c  sw $s0,80($zero)
        32:     data <= 32'h20100003;    //0x80  addi $s0,$zero,3
        33:     data <= 32'hac100054;    //0x84  sw $s0,84($zero)
        34:     data <= 32'h20100046;    //0x88  addi $s0,$zero,70
        35:     data <= 32'hac100058;    //0x8c  sw $s0,88($zero)
        36:     data <= 32'h20100021;    //0x90  addi $s0,$zero,33
        37:     data <= 32'hac10005c;    //0x94  sw $s0,92($zero)
        38:     data <= 32'h20100006;    //0x98  addi $s0,$zero,6
        39:     data <= 32'hac100060;    //0x9c  sw $s0,96($zero)
        40:     data <= 32'h2010000e;    //0xa0  addi $s0,$zero,14
        41:     data <= 32'hac100064;    //0xa4  sw $s0,100($zero)
        42:     data <= 32'h20030001;    //0xa8  addi $v1,$zero,1
        43:     data <= 32'h08000077;    //0xac  j End
        44:     data <= 32'h20080003;    //0xb0  addi $t0,$zero,3
        45:     data <= 32'haec80008;    //0xb4  sw $t0,8($s6)
        46:     data <= 32'h00035842;    //0xb8  srl $t3,$v1,1
        47:     data <= 32'h11600006;    //0xbc  beq $t3,$zero,A
        48:     data <= 32'h000b5842;    //0xc0  srl $t3,$t3,1
        49:     data <= 32'h1160000d;    //0xc4  beq $t3,$zero,B
        50:     data <= 32'h000b5842;    //0xc8  srl $t3,$t3,1
        51:     data <= 32'h11600014;    //0xcc  beq $t3,$zero,C
        52:     data <= 32'h000b5842;    //0xd0  srl $t3,$t3,1
        53:     data <= 32'h1160001b;    //0xd4  beq $t3,$zero,D
        54:     data <= 32'h8ecc0018;    //0xd8  lw $t4,24($s6)
        55:     data <= 32'h318c000f;    //0xdc  andi $t4,$t4,15
        56:     data <= 32'h000c6080;    //0xe0  sll $t4,$t4,2
        57:     data <= 32'h8d8c0028;    //0xe4  lw $t4,40($t4)
        58:     data <= 32'h00036a00;    //0xe8  sll $t5,$v1,8
        59:     data <= 32'h01ac6020;    //0xec  add $t4,$t5,$t4
        60:     data <= 32'haecc0014;    //0xf0  sw $t4,20($s6)
        61:     data <= 32'h20030002;    //0xf4  addi $v1,$zero,2
        62:     data <= 32'h0800005a;    //0xf8  j cycle
        63:     data <= 32'h8ecc0018;    //0xfc  lw $t4,24($s6)
        64:     data <= 32'h318c00f0;    //0x100 andi $t4,$t4,240
        65:     data <= 32'h000c6082;    //0x104 srl $t4,$t4,2
        66:     data <= 32'h8d8c0028;    //0x108 lw $t4,40($t4)
        67:     data <= 32'h00036a00;    //0x10c sll $t5,$v1,8
        68:     data <= 32'h01ac6020;    //0x110 add $t4,$t5,$t4
        69:     data <= 32'haecc0014;    //0x114 sw $t4,20($s6)
        70:     data <= 32'h20030004;    //0x118 addi $v1,$zero,4
        71:     data <= 32'h0800005a;    //0x11c j cycle
        72:     data <= 32'h8ecc001c;    //0x120 lw $t4,28($s6)
        73:     data <= 32'h318c000f;    //0x124 andi $t4,$t4,15
        74:     data <= 32'h000c6080;    //0x128 sll $t4,$t4,2
        75:     data <= 32'h8d8c0028;    //0x12c lw $t4,40($t4)
        76:     data <= 32'h00036a00;    //0x130 sll $t5,$v1,8
        77:     data <= 32'h01ac6020;    //0x134 add $t4,$t5,$t4
        78:     data <= 32'haecc0014;    //0x138 sw $t4,20($s6)
        79:     data <= 32'h20030008;    //0x13c addi $v1,$zero,8
        80:     data <= 32'h0800005a;    //0x140 j cycle
        81:     data <= 32'h8ecc001c;    //0x144 lw $t4,28($s6)
        82:     data <= 32'h318c00f0;    //0x148 andi $t4,$t4,240
        83:     data <= 32'h000c6082;    //0x14c srl $t4,$t4,2
        84:     data <= 32'h8d8c0028;    //0x150 lw $t4,40($t4)
        85:     data <= 32'h00036a00;    //0x154 sll $t5,$v1,8
        86:     data <= 32'h01ac6020;    //0x158 add $t4,$t5,$t4
        87:     data <= 32'haecc0014;    //0x15c sw $t4,20($s6)
        88:     data <= 32'h20030001;    //0x160 addi $v1,$zero,1
        89:     data <= 32'h0800005a;    //0x164 j cycle
        90:     data <= 32'h8ec80024;    //0x168 lw $t0,36($s6)
        91:     data <= 32'h000847c0;    //0x16c sll $t0,$t0,31
        92:     data <= 32'h000847c2;    //0x170 srl $t0,$t0,31
        93:     data <= 32'h11000017;    //0x174 beq $t0,$zero,InEnd
        94:     data <= 32'h00004020;    //0x178 add $t0,$zero,$zero
        95:     data <= 32'haec80024;    //0x17c sw $t0,36($s6)
        96:     data <= 32'h8ec90018;    //0x180 lw $t1,24($s6)
        97:     data <= 32'h8eca001c;    //0x184 lw $t2,28($s6)
        98:     data <= 32'h11200008;    //0x188 beq $t1,$zero,end1
        99:     data <= 32'h11400007;    //0x18c beq $t2,$zero,end1
        100:    data <= 32'h112a0007;    //0x190 beq $t1,$t2,end2
        101:    data <= 32'h0149402a;    //0x194 slt $t0,$t2,$t1
        102:    data <= 32'h11000002;    //0x198 beq $t0,$zero,loop2
        103:    data <= 32'h012a4822;    //0x19c sub $t1,$t1,$t2
        104:    data <= 32'h08000064;    //0x1a0 j loop1
        105:    data <= 32'h01495022;    //0x1a4 sub $t2,$t2,$t1
        106:    data <= 32'h08000064;    //0x1a8 j loop1
        107:    data <= 32'h00005020;    //0x1ac add $t2,$zero,$zero
        108:    data <= 32'h01401020;    //0x1b0 add $v0,$t2,$zero
        109:    data <= 32'haec20020;    //0x1b4 sw $v0,32($s6)
        110:    data <= 32'haec2000c;    //0x1b8 sw $v0,12($s6)
        111:    data <= 32'h8ec80024;    //0x1bc lw $t0,36($s6)
        112:    data <= 32'h00084082;    //0x1c0 srl $t0,$t0,2
        113:    data <= 32'h15000003;    //0x1c4 bne $t0,$zero,InEnd
        114:    data <= 32'h200a0002;    //0x1c8 addi $t2,$zero,2
        115:    data <= 32'haeca0024;    //0x1cc sw $t2,36($s6)
        116:    data <= 32'h00000000;    //0x1d0 sll $zero,$zero,0
        117:    data <= 32'h03400008;    //0x1d4 jr $k0
        118:    data <= 32'h03400008;    //0x1d8 jr $k0
        119:    data <= 32'h08000077;    //0x1dc j End
      default:  data <= 32'h08000000;
    endcase
endmodule
